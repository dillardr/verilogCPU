`include "parameter.v"

//enables 32 registers

//rs = register select
//ws = write select
//wd =
//rd = register d
//we =

module gpreg(
    input[]

)