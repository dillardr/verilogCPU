`include "parameter.v"

module instreg(
    input[`col-1:0] addr,
    output[`col-1:0] inst

);


//Sets up memory and loads instruction from file


endmodule