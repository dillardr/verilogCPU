`include "parameter.v"

module datamemory (
    input[`col -1:0] addr, data_in,
    input clk,
    input we,
    output[`col -1: 0] data
);
    
endmodule