
module adder(
    output reg[15:0] out,
    input [7:0] ina, inb,
    input clk, sclrn

);




endmodule 
