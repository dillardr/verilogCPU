`include "parameter.v"


module instreg(
    input [`col-1:0] inst_in,
    output [`col-1:0] inst_out
);

endmodule