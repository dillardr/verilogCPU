`include "parameter.v"

module instdecode (
    input [`col-1:0] inst_in,
    input clk,
    //outputs will be added as funtions are added
);
    
endmodule

