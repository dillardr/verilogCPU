`include "parameter.v"

module progcount (
    input [`col-1:0] count_in,
    input clk, we,
    output [`col-1:0] count_out,
);
    
endmodule